module xor_gate (A,B,y);
    input A,B;
    output y;
   xor(y,A,B);
endmodule