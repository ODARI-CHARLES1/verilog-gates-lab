module and_gate (A,B,y);
    input A,B;
    output y;
    and(y,A,B);
endmodule