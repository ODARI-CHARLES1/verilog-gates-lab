module not_gate (A,y);
    input A;
    output y;
    not(y,A);
endmodule