module xnor_gate (A,B,y);
    input A,B;
    output y;
    xnor(y,A,B);
endmodule