
module nand_gate (A,B,y);
    input A,B;
    output y;
    nand(y,A,B);
endmodule